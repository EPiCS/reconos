library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity invSbox is
	port(
	  clk       : in std_logic;
	  rst       : in std_logic;
		addr      : in	STD_LOGIC_VECTOR  (7 downto 0);	  -- Byte
		sByte     : out STD_LOGIC_VECTOR (7 downto 0)	 -- Substituted Byte		
		);		
end invSbox;


architecture invSbox of invSbox is
TYPE byte_array is array(0 to 255) of std_logic_vector (7 downto 0);
constant memory: byte_array:=(
		0	=> X"52", 1 => X"09", 2 => X"6A", 3 => X"D5", 4 => X"30", 5 => X"36", 6 => X"A5", 7 => X"38",
		8	=> X"BF", 9 => X"40", 10 => X"A3", 11 => X"9E", 12 => X"81", 13 => X"F3", 14 => X"D7", 15 => X"FB",
		16	=> X"7C", 17 => X"E3", 18 => X"39", 19 => X"82", 20 => X"9B", 21 => X"2F", 22 => X"FF", 23 => X"87",
		24	=> X"34", 25 => X"8E", 26 => X"43", 27 => X"44", 28 => X"C4", 29 => X"DE", 30 => X"E9", 31 => X"CB",
		32	=> X"54", 33 => X"7B", 34 => X"94", 35 => X"32", 36 => X"A6", 37 => X"C2", 38 => X"23", 39 => X"3D",
		40	=> X"EE", 41 => X"4C", 42 => X"95", 43 => X"0B", 44 => X"42", 45 => X"FA", 46 => X"C3", 47 => X"4E",
		48	=> X"08", 49 => X"2E", 50 => X"A1", 51 => X"66", 52 => X"28", 53 => X"D9", 54 => X"24", 55 => X"B2",
		56	=> X"76", 57 => X"5B", 58 => X"A2", 59 => X"49", 60 => X"6D", 61 => X"8B", 62 => X"D1", 63 => X"25",
		64	=> X"72", 65 => X"F8", 66 => X"F6", 67 => X"64", 68 => X"86", 69 => X"68", 70 => X"98", 71 => X"16",
		72	=> X"D4", 73 => X"A4", 74 => X"5C", 75 => X"CC", 76 => X"5D", 77 => X"65", 78 => X"B6", 79 => X"92",
		80	=> X"6C", 81 => X"70", 82 => X"48", 83 => X"50", 84 => X"FD", 85 => X"ED", 86 => X"B9", 87 => X"DA",
		88	=> X"5E", 89 => X"15", 90 => X"46", 91 => X"57", 92 => X"A7", 93 => X"8D", 94 => X"9D", 95 => X"84",
		96	=> X"90", 97 => X"D8", 98 => X"AB", 99 => X"00", 100 => X"8C", 101 => X"BC", 102 => X"D3", 103 => X"0A",
		104 => X"F7", 105 => X"E4", 106 => X"58", 107 => X"05", 108 => X"B8", 109 => X"B3", 110 => X"45", 111 => X"06",
		112 => X"D0", 113 => X"2C", 114 => X"1E", 115 => X"8F", 116 => X"CA", 117 => X"3F", 118 => X"0F", 119 => X"02",
		120 => X"C1", 121 => X"AF", 122 => X"BD", 123 => X"03", 124 => X"01", 125 => X"13", 126 => X"8A", 127 => X"6B",
		128 => X"3A", 129 => X"91", 130 => X"11", 131 => X"41", 132 => X"4F", 133 => X"67", 134 => X"DC", 135 => X"EA",
		136 => X"97", 137 => X"F2", 138 => X"CF", 139 => X"CE", 140 => X"F0", 141 => X"B4", 142 => X"E6", 143 => X"73",
		144 => X"96", 145 => X"AC", 146 => X"74", 147 => X"22", 148 => X"E7", 149 => X"AD", 150 => X"35", 151 => X"85",
		152 => X"E2", 153 => X"F9", 154 => X"37", 155 => X"E8", 156 => X"1C", 157 => X"75", 158 => X"DF", 159 => X"6E",
		160 => X"47", 161 => X"F1", 162 => X"1A", 163 => X"71", 164 => X"1D", 165 => X"29", 166 => X"C5", 167 => X"89",
		168 => X"6F", 169 => X"B7", 170 => X"62", 171 => X"0E", 172 => X"AA", 173 => X"18", 174 => X"BE", 175 => X"1B",
		176 => X"FC", 177 => X"56", 178 => X"3E", 179 => X"4B", 180 => X"C6", 181 => X"D2", 182 => X"79", 183 => X"20",
		184 => X"9A", 185 => X"DB", 186 => X"C0", 187 => X"FE", 188 => X"78", 189 => X"CD", 190 => X"5A", 191 => X"F4",
		192 => X"1F", 193 => X"DD", 194 => X"A8", 195 => X"33", 196 => X"88", 197 => X"07", 198 => X"C7", 199 => X"31",
		200 => X"B1", 201 => X"12", 202 => X"10", 203 => X"59", 204 => X"27", 205 => X"80", 206 => X"EC", 207 => X"5F",
		208 => X"60", 209 => X"51", 210 => X"7F", 211 => X"A9", 212 => X"19", 213 => X"B5", 214 => X"4A", 215 => X"0D",
		216 => X"2D", 217 => X"E5", 218 => X"7A", 219 => X"9F", 220 => X"93", 221 => X"C9", 222 => X"9C", 223 => X"EF",
		224 => X"A0", 225 => X"E0", 226 => X"3B", 227 => X"4D", 228 => X"AE", 229 => X"2A", 230 => X"F5", 231 => X"B0",
		232 => X"C8", 233 => X"EB", 234 => X"BB", 235 => X"3C", 236 => X"83", 237 => X"53", 238 => X"99", 239 => X"61",
		240 => X"17", 241 => X"2B", 242 => X"04", 243 => X"7E", 244 => X"BA", 245 => X"77", 246 => X"D6", 247 => X"26",
		248 => X"E1", 249 => X"69", 250 => X"14", 251 => X"63", 252 => X"55", 253 => X"21", 254 => X"0C", 255 => X"7D"
		);

begin

process(rst, addr)
  begin
    if(rst='1')then
      sByte<=X"00";
    else
      sByte<=memory(to_integer(unsigned(addr)));
    end if;
end process;
      
end invSbox;
