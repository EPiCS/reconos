../../ise_project/system/system_top.vhd