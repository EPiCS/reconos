

-- @module : shadowing_control
-- @author : meise
-- @date   : 23.05.2016


library ieee;
use ieee.std_logic_1164.all;

entity shadowing_control is 
port (
    clk			: in	  std_logic); 
     
end shadowing_control;     
        

architecture synth of shadowing_control is
               
begin  

-- control muxes and sh_units and relay error messages

end synth;








