/home/meise/git/reconos_epics/externals/easics/PCK_CRC32_D32.vhd